    module level_one (
        input  logic [5:0] addr,
        output logic [39:0] data
    );
    // 30 rows, 40 columns
        always_comb begin
            case (addr)
                6'd0:  data = 40'b0000000000000000000000000000000000000000;
                6'd1:  data = 40'b0000000000000000000000000000000000000000;
                6'd2:  data = 40'b0000000001111100001111100111110000000000;
                6'd3:  data = 40'b0000000001111100011111100111110000000000;
                6'd4:  data = 40'b0000000001100000011100000110000000000000;
                6'd5:  data = 40'b0000000001100000011000000110000000000000;
                6'd6:  data = 40'b0000000001111000011000000111100000000000;
                6'd7:  data = 40'b0000000001111000011000000111100000000000;
                6'd8:  data = 40'b0000000001100000011000000110000000000000;
                6'd9:  data = 40'b0000000001100000011100000110000000000000;
                6'd10: data = 40'b0000000001111100011111100111110000000000;
                6'd11: data = 40'b0000000001111100001111100111110000000000;
                6'd12: data = 40'b0000000000000000000000000000000000000000;
                6'd13: data = 40'b0000000000000000000000000000000000000000;
                6'd14: data = 40'b0000000111110000011111100001111110000000;
                6'd15: data = 40'b0000000111110000011001100001111110000000;
                6'd16: data = 40'b0000000000110000011001100001100000000000;
                6'd17: data = 40'b0000000000110000011001100001100000000000;
                6'd18: data = 40'b0000000111110000011111100001111110000000;
                6'd19: data = 40'b0000000111110000011111100001111110000000;
                6'd20: data = 40'b0000000000110000011001100000000110000000;
                6'd21: data = 40'b0000000000110000011001100000000110000000;
                6'd22: data = 40'b0000000111110000011001100001111110000000;
                6'd23: data = 40'b0000000111110000011111100001111110000000;
                6'd24: data = 40'b0000000000000000000000000000000000000000;
                6'd25: data = 40'b0000000000000000000000000000000000000000;
                6'd26: data = 40'b0000000000000000000000000000000000000000;
                6'd27: data = 40'b0000000000000000001111000000000000000000;
                6'd28: data = 40'b0000000000000000001001000000000000000000;
                6'd29: data = 40'b0000000000000000001001000000000000000000;
                default: data = 40'b0;
            endcase
        end
    endmodule

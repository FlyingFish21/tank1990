module heart_example (
	input logic vga_clk,
	input logic [9:0] DrawX, DrawY,
	input logic show_heart,
	output logic [3:0] red, green, blue
);

logic [6:0] rom_address;
logic [1:0] rom_q;

logic [3:0] palette_red, palette_green, palette_blue;

logic negedge_vga_clk;

// read from ROM on negedge, set pixel on posedge
assign negedge_vga_clk = ~vga_clk;

// address into the rom = (x*xDim)/640 + ((y*yDim)/480) * xDim
// this will stretch out the sprite across the entire screen
assign rom_address = ((DrawX * 11) / 640) + (((DrawY * 11) / 480) * 11);

always_ff @ (posedge vga_clk) begin
	red <= 4'h0;
	green <= 4'h0;
	blue <= 4'h0;

	if (show_heart) begin
		red <= palette_red;
		green <= palette_green;
		blue <= palette_blue;
	end
end

heart_rom heart_rom (
	.clka   (negedge_vga_clk),
	.addra (rom_address),
	.douta       (rom_q)
);

heart_palette heart_palette (
	.index (rom_q),
	.red   (palette_red),
	.green (palette_green),
	.blue  (palette_blue)
);

endmodule
